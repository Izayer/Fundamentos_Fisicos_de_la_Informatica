* Carga condensadores
v0 0 1 type=vdc vdc=10
r1 3 1 3k
c1 0 2 47u ic=0
v1dummy 2 3 type=vdc vdc=0
c2 0 4 22u ic=0
v2dummy 4 3 type=vdc vdc=0
.op
.tran tstep=0.01 tstop=1 uic=0
.end
